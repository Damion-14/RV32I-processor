module alu_ctl(
  input wire [ 5:0 ] alu_op,
  input wire [ 31:0 ] instruction,

  output wire [ 2:0 ] i_opsel,
  output wire i_sub, 
  output wire i_unsigned, 
  output wire i_arith,

);
// TODO 

endmodule